module test (
    input a,
    output [1:0] b
    );

assign a = b + 1;

endmodule
