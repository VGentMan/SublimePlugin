 wad <= -234